module top_key_led(
    input      wire sys_clk,
    input      wire sys_rst_n,
    input      wire key_in_raw,     // ��Ӧ������KEY1
    output     reg  led_out         //��Ӧled
);

    wire key_pressed_pulse;//������������ź�
    
    //ʵ��������ģ��
    
    key_debounce u_debounce(
        .sys_clk    (sys_clk),
        .sys_rst_n  (sys_rst_n),
        .key_in     (key_in_raw),
        .key_flag   (key_pressed_pulse),//���������ź�
        .key_value  ()
    );
    
    always @(posedge sys_clk or negedge sys_rst_n)begin
        if(!sys_rst_n)begin
            led_out <= 1'b1;
        end 
        else if(key_pressed_pulse)begin
            led_out <= ~led_out; 
        end
    end
    
endmodule

        