module div_3(
    input           clk_in,
    input           rst_n,
    output          clk_out
);

    reg [1:0] r_cnt;

    // 1. �������߼� (������ԭ����д��)
    always @(posedge clk_in or negedge rst_n) begin
        if(!rst_n)
            r_cnt <= 2'd0;
        else 
            r_cnt <= (r_cnt == 2'd2) ? 2'd0 : r_cnt + 1;
    end

    reg clk_p;
    reg clk_n;

    // 2. �����ز������� clk_p
    // ������Ϊ 2 ʱ���ߣ�����ʱ������ (�ߵ�ƽռ 1/3)
    always @(posedge clk_in or negedge rst_n) begin
        if(!rst_n)
            clk_p <= 1'b0;
        else if (r_cnt == 2'd2) 
            clk_p <= 1'b1;
        else 
            clk_p <= 1'b0;
    end

    // 3. �½��ز������� clk_n
    // ͬ���ڼ���Ϊ 2 ʱ���� (ע�⣺r_cnt ���������ر�ģ��������½��ز����� r_cnt ֵ���� 2)
    always @(negedge clk_in or negedge rst_n) begin
        if(!rst_n)
            clk_n <= 1'b0;
        else if (r_cnt == 2'd2) 
            clk_n <= 1'b1;
        else 
            clk_n <= 1'b0;
    end

    // 4. ������
    // ��������ڵ����������ࡰ�򡱣��õ� 1.5 �����ڵĸߵ�ƽ
    assign clk_out = clk_p | clk_n;

endmodule

// generate testbench for module div_3
