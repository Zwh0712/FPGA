module seg_driver(
    input             sys_clk,      
    input             sys_rst_n,    
    input      [15:0] data_in,      
    input      [3:0]  point_on,     
    output reg [3:0]  seg_sel,      
    output reg [7:0]  seg_led       
);

    parameter CNT_MAX = 16'd49_999; 

    // 1. ɨ�趨ʱ�� (����)
    reg [15:0] cnt_scan;
    wire       scan_tick;
    always @(posedge sys_clk or negedge sys_rst_n) begin
        if (!sys_rst_n) cnt_scan <= 16'd0;
        else if (cnt_scan == CNT_MAX) cnt_scan <= 16'd0;
        else cnt_scan <= cnt_scan + 1'b1;
    end
    assign scan_tick = (cnt_scan == CNT_MAX);

    // 2. ״̬�л� (����)
    reg [1:0] state; 
    always @(posedge sys_clk or negedge sys_rst_n) begin
        if (!sys_rst_n) state <= 2'd0;
        else if (scan_tick) state <= state + 1'b1;
    end

    // 3. λѡ�߼� (*** �޸ĵ� 1����Ϊ�������߼� ***)
    // �������������˽ӵ�(0)Ϊѡ�У���ѡ�и�(1)
    
    reg [3:0] num_disp; 
    reg       dot_disp; 

    always @(*) begin
        case (state)
            2'd0: begin 
                seg_sel  = 4'b1110;          // <--- �޸ģ�0ѡ�е�0λ
                num_disp = data_in[3:0];     
                dot_disp = point_on[0];      
            end
            2'd1: begin 
                seg_sel  = 4'b1101;          // <--- �޸ģ�0ѡ�е�1λ
                num_disp = data_in[7:4];
                dot_disp = point_on[1];
            end
            2'd2: begin 
                seg_sel  = 4'b1011;          // <--- �޸ģ�0ѡ�е�2λ
                num_disp = data_in[11:8];
                dot_disp = point_on[2];
            end
            2'd3: begin 
                seg_sel  = 4'b0111;          // <--- �޸ģ�0ѡ�е�3λ
                num_disp = data_in[15:12];
                dot_disp = point_on[3];
            end
            default: begin
                seg_sel  = 4'b1111;          // ȫ��ѡ
                num_disp = 4'd0;
                dot_disp = 1'b0;
            end
        endcase
    end

    // 4. �������� (���䣬���ζ��屾���Ǹߵ�ƽ��Ч��)
    reg [6:0] seg_decode; 
    always @(*) begin
        case (num_disp)
            4'h0: seg_decode = 7'b011_1111; 
            4'h1: seg_decode = 7'b000_0110; 
            4'h2: seg_decode = 7'b101_1011; 
            4'h3: seg_decode = 7'b100_1111; 
            4'h4: seg_decode = 7'b110_0110; 
            4'h5: seg_decode = 7'b110_1101; 
            4'h6: seg_decode = 7'b111_1101; 
            4'h7: seg_decode = 7'b000_0111; 
            4'h8: seg_decode = 7'b111_1111; 
            4'h9: seg_decode = 7'b110_1111; 
            4'hA: seg_decode = 7'b111_0111; 
            4'hB: seg_decode = 7'b111_1100; 
            4'hC: seg_decode = 7'b011_1001; 
            4'hD: seg_decode = 7'b101_1110; 
            4'hE: seg_decode = 7'b111_1001; 
            4'hF: seg_decode = 7'b111_0001; 
            default: seg_decode = 7'b000_0000;
        endcase
    end

    // 5. �������ƴװ (*** �޸ĵ� 2������������Ҫȡ�� ***)
    // ����������ѡ���ߵ�ƽ(1)����
    always @(*) begin
        // ȥ���˲��˺� ~
        seg_led = {dot_disp, seg_decode}; 
    end

endmodule
