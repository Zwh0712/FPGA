module led_multi_clock(
    input  wire sys_clk,      // ϵͳʱ�� 50MHz
    input  wire sys_rst_n,    // ϵͳ��λ (�͵�ƽ��Ч)
    output reg  [1:0] led     // 2��LED��
);

    // ����ʱ�䳣�� (50MHzʱ����)
    // 0.5�� = 25,000,000 ������
    parameter CNT_MAX_0 = 26'd24_999_999; 
    // 0.25�� = 12,500,000 ������
    parameter CNT_MAX_1 = 26'd12_499_999;

    // ��������������
    reg [25:0] cnt0;
    reg [25:0] cnt1;

    // ---------------------------------------------------------
    // �߼���1������ LED[0] (����: 0.5s ��ת)
    // ---------------------------------------------------------
    always @(posedge sys_clk or negedge sys_rst_n) begin
        if (!sys_rst_n) begin
            cnt0   <= 26'd0;
            led[0] <= 1'b1;  // ��λʱ�� (����ߵ�ƽ�����ӵ�·������ͨ��ZYNQ���Ǹߵ�ƽ��)
        end
        else if (cnt0 == CNT_MAX_0) begin
            cnt0   <= 26'd0;
            led[0] <= ~led[0]; // ��ת״̬
        end
        else begin
            cnt0   <= cnt0 + 1'b1;
        end
    end

    // ---------------------------------------------------------
    // �߼���2������ LED[1] (����: 0.25s ��ת)
    // ---------------------------------------------------------
    always @(posedge sys_clk or negedge sys_rst_n) begin
        if (!sys_rst_n) begin
            cnt1   <= 26'd0;
            led[1] <= 1'b0;  // ��λʱ�� (�������ó�ʼ״̬��ͬ)
        end
        else if (cnt1 == CNT_MAX_1) begin
            cnt1   <= 26'd0;
            led[1] <= ~led[1]; // ��ת״̬
        end
        else begin
            cnt1   <= cnt1 + 1'b1;
        end
    end

endmodule