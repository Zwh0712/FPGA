module key_debounce(
    input   wire  sys_clk,      //50MHz
    input   wire  sys_rst_n,
    input   wire  key_in,       //���������루���ܴ�������
    
    output  reg  key_flag,   //�����һ��ʱ�����ڵ����壬��������Ч����
    output  reg  key_value   //�������������ȶ���ƽ
);

    //20ms ������Ŀ��ֵ
    //50MHz *0.02s = 1000000
    parameter CNT_MAX = 20'd1_000_000;
    
    reg [19:0] cnt;
    reg key_reg;
    
    //״̬��/�������߼�
    always@(posedge sys_clk or negedge sys_rst_n) begin
        if(!sys_rst_n)begin
            cnt       <= 20'd0;
            key_flag  <= 1'b0;
            key_value <= 1'b1;  //Ĭ�ϸߵ�ƽ��δ���£�
        end
        else begin
        //Ĭ�Ͻ���־λ���ͣ�ֻ���ڼ�������һ˲������
        key_flag      <= 1'b0;
        //��������ǵ͵�ƽ�����谴��Ϊ0��
        if(key_in == 1'b0)begin
            //�����������û������һֱ��
            if(cnt < CNT_MAX)begin
                cnt <= cnt + 1'b1;
            end
            //�պ�����20ms ����һ��
            else if (cnt == CNT_MAX)begin
                key_flag    <= 1'b1;
                key_value   <= 1'b0;
                cnt         <= cnt + 1'b1;
            end
            //  �������󣬱�����״��ʲô��������ֱ���ɿ�����
        end
        else begin
            //  ����һ����ߣ��ɿ��򶶶�����ߣ����������������㣡
            //  ����ǡ��������ĺ��ģ����������͵�ƽ���м��һ�¾�Ҫ������
            cnt          <= 20'd0;
            key_value    <= 1'b1;
        end
    end
end

endmodule

        
            